wire [3 : 0]  m_axi_awid    ;
wire [30 : 0] m_axi_awaddr  ;
wire [7 : 0]  m_axi_awlen   ;
wire [2 : 0]  m_axi_awsize  ;
wire [1 : 0]  m_axi_awburst ;
wire [0 : 0]  m_axi_awlock  ;
wire [3 : 0]  m_axi_awcache ;
wire [2 : 0]  m_axi_awprot  ;
wire [3 : 0]  m_axi_awqos   ;
wire [3 : 0]  m_axi_awregion;
wire          m_axi_awvalid ;
wire          m_axi_awready ;
wire [63 : 0] m_axi_wdata   ;
wire [7 : 0]  m_axi_wstrb   ;
wire          m_axi_wlast   ;
wire          m_axi_wvalid  ;
wire          m_axi_wready  ;
wire [3 : 0]  m_axi_bid     ;
wire [1 : 0]  m_axi_bresp   ;
wire          m_axi_bvalid  ;
wire          m_axi_bready  ;
wire [3 : 0]  m_axi_arid    ;
wire [30 : 0] m_axi_araddr  ;
wire [7 : 0]  m_axi_arlen   ;
wire [2 : 0]  m_axi_arsize  ;
wire [1 : 0]  m_axi_arburst ;
wire [0 : 0]  m_axi_arlock  ;
wire [3 : 0]  m_axi_arcache ;
wire [2 : 0]  m_axi_arprot  ;
wire [3 : 0]  m_axi_arqos   ;
wire [3 : 0]  m_axi_arregion;
wire          m_axi_arvalid ;
wire          m_axi_arready ;
wire [3 : 0]  m_axi_rid     ;
wire [63 : 0] m_axi_rdata   ;
wire [1 : 0]  m_axi_rresp   ;
wire          m_axi_rlast   ;
wire          m_axi_rvalid  ;
wire          m_axi_rready  ;