input  wire[19 : 0] s_axi_awaddr,
input  wire[7 : 0]  s_axi_awlen,
input  wire[2 : 0]  s_axi_awsize,
input  wire[1 : 0]  s_axi_awburst,
input  wire         s_axi_awlock,
input  wire[3 : 0]  s_axi_awcache,
input  wire[2 : 0]  s_axi_awprot,
input  wire         s_axi_awvalid,
output wire         s_axi_awready,
input  wire[31 : 0] s_axi_wdata,
input  wire[3 : 0]  s_axi_wstrb,
input  wire         s_axi_wlast,
input  wire         s_axi_wvalid,
output wire         s_axi_wready,
output wire[1 : 0]  s_axi_bresp,
output wire         s_axi_bvalid,
input  wire         s_axi_bready,
input  wire[19 : 0] s_axi_araddr,
input  wire[7 : 0]  s_axi_arlen,
input  wire[2 : 0]  s_axi_arsize,
input  wire[1 : 0]  s_axi_arburst,
input  wire         s_axi_arlock,
input  wire[3 : 0]  s_axi_arcache,
input  wire[2 : 0]  s_axi_arprot,
input  wire         s_axi_arvalid,
output wire         s_axi_arready,
output wire[31 : 0] s_axi_rdata,
output wire[1 : 0]  s_axi_rresp,
output wire         s_axi_rlast,
output wire         s_axi_rvalid,
input  wire         s_axi_rready