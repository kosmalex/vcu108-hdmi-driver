.s_axi_awaddr  (m_axi_awaddr ),
.s_axi_awlen   (m_axi_awlen  ),
.s_axi_awsize  (m_axi_awsize ),
.s_axi_awburst (m_axi_awburst),
.s_axi_awlock  (m_axi_awlock ),
.s_axi_awcache (m_axi_awcache),
.s_axi_awprot  (m_axi_awprot ),
.s_axi_awvalid (m_axi_awvalid),
.s_axi_awready (m_axi_awready),
.s_axi_wdata   (m_axi_wdata  ),
.s_axi_wstrb   (m_axi_wstrb  ),
.s_axi_wlast   (m_axi_wlast  ),
.s_axi_wvalid  (m_axi_wvalid ),
.s_axi_wready  (m_axi_wready ),
.s_axi_bresp   (m_axi_bresp  ),
.s_axi_bvalid  (m_axi_bvalid ),
.s_axi_bready  (m_axi_bready ),

.s_axi_araddr  ('d0 ),
.s_axi_arlen   ('d0 ),
.s_axi_arsize  ('d0 ),
.s_axi_arburst ('d0 ),
.s_axi_arlock  ('d0 ),
.s_axi_arcache ('d0 ),
.s_axi_arprot  ('d0 ),
.s_axi_arvalid (1'b0),
.s_axi_arready (    ),
.s_axi_rdata   (    ),
.s_axi_rresp   (    ),
.s_axi_rlast   (    ),
.s_axi_rvalid  (    ),
.s_axi_rready  (1'b0),