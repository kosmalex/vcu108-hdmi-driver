logic[31 : 0] m_axi_awaddr  ;
logic[7 : 0]  m_axi_awlen   ;
logic[2 : 0]  m_axi_awsize  ;
logic[1 : 0]  m_axi_awburst ;
logic[0 : 0]  m_axi_awlock  ;
logic[3 : 0]  m_axi_awcache ;
logic[2 : 0]  m_axi_awprot  ;
logic[3 : 0]  m_axi_awqos   ;
logic[3 : 0]  m_axi_awregion;
logic         m_axi_awvalid ;
logic         m_axi_awready ;
logic[31 : 0] m_axi_wdata   ;
logic[3 : 0]  m_axi_wstrb   ;
logic         m_axi_wlast   ;
logic         m_axi_wvalid  ;
logic         m_axi_wready  ;
logic[1 : 0]  m_axi_bresp   ;
logic         m_axi_bvalid  ;
logic         m_axi_bready  ;